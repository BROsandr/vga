// The module converts axil input interface to simple native out interface.

module vga_axil_slave_fsm
  import vga_axil_pkg::axil_data_t, vga_axil_pkg::axil_addr_t, vga_axil_pkg::native_addr_t;
(
  vga_axil_if.slave axil_if,
  vga_native_if     native_if
);

// START fsm state_ff, state_next logic
  localparam int  NUM_OF_STATES = 5;
  localparam type state_e = enum bit [$clog2(NUM_OF_STATES)-1:0] {
    StIdle,
    StAddr,
    StData,
    StResp,
    StAddrData
  };
  state_e read_state_ff, read_state_next, write_state_ff, write_state_next;

  always_ff @(posedge axil_if.clk_i or negedge axil_if.arst_ni) begin
    if (!axil_if.arst_ni) begin
      read_state_ff  <= StIdle;
      write_state_ff <= StIdle;
    end else begin
      read_state_ff  <= read_state_next;
      write_state_ff <= write_state_next;
    end
  end

  // state_ff is indicating what has already been done.
  //   For example state == StAddr indicates that an address has been accepted.
  always_comb begin : read
    read_state_next = read_state_ff;
    unique case (read_state_ff)
      StIdle: if (axil_if.ar_handshake_i) read_state_next = StAddr;
      StAddr:                             read_state_next = StData;
      StData:                             read_state_next = StResp;
      StResp: if (axil_if.r_handshake_i)  read_state_next = StIdle;

      default:                            read_state_next = StIdle;
    endcase
  end

  always_comb begin : write
    write_state_next = write_state_ff;
    unique case (write_state_ff)
      StIdle    : if (axil_if.aw_handshake_i && axil_if.w_handshake_i) write_state_next = StAddrData;
      StAddrData:                                                      write_state_next = StResp;
      StResp    : if (axil_if.b_handshake_i)                           write_state_next = StIdle;

      default:                                                         write_state_next = StIdle;
    endcase
  end
// END fsm state_ff, state_next logic

// START read logic
// START axil_if.arready
  logic arready_ff;
  logic arready_next;

  assign arready_next = read_state_next == StIdle;

  always_ff @(posedge axil_if.clk_i or negedge axil_if.arst_ni) begin
    if      (!axil_if.arst_ni) arready_ff <= '0;
    else                       arready_ff <= arready_next;
  end
// END axil_if.arready

// START addr_read_ff
  native_addr_t addr_read_ff;
  native_addr_t addr_read_next;
  logic         addr_read_en;

  assign      addr_read_en   = read_state_next == StAddr;

  import      vga_axil_pkg::axil2native_addr;
  assign      addr_read_next = axil2native_addr(axil_if.araddr_i);

  always_ff @(posedge axil_if.clk_i or negedge axil_if.arst_ni) begin
    if      (!axil_if.arst_ni) addr_read_ff <= '0;
    else if (addr_read_en    ) addr_read_ff <= addr_read_next;
  end
// END addr_read_ff

// START read_en_sync
  logic read_en_sync_ff;
  logic read_en_sync_next;

  assign read_en_sync_next = read_state_next == StAddr;

  always_ff @(posedge axil_if.clk_i or negedge axil_if.arst_ni) begin
    if      (!axil_if.arst_ni) read_en_sync_ff <= '0;
    else                       read_en_sync_ff <= read_en_sync_next;
  end
// END read_en_sync

// START axil_if.rrvalid
  logic rvalid_ff;
  logic rvalid_next;

  assign rvalid_next = read_state_next == StResp;

  always_ff @(posedge axil_if.clk_i or negedge axil_if.arst_ni) begin
    if      (!axil_if.arst_ni) rvalid_ff <= '0;
    else                       rvalid_ff <= rvalid_next;
  end
// END axil_if.rvalid

// START axil_if.rdata
  axil_data_t rdata_ff;
  axil_data_t rdata_next;
  logic       rdata_en;

  assign rdata_en   = read_state_next == StResp;
  assign rdata_next = native_if.data2axil;

  always_ff @(posedge axil_if.clk_i or negedge axil_if.arst_ni) begin
    if      (!axil_if.arst_ni) rdata_ff <= '0;
    else if (rdata_en        ) rdata_ff <= rdata_next;
  end
// END axil_if.rdata
// END read logic

// START write logic
// START write_en
  logic write_en_ff;
  logic write_en_next;

  assign write_en_next = write_state_next == StAddrData;

  always_ff @(posedge axil_if.clk_i or negedge axil_if.arst_ni) begin
    if      (!axil_if.arst_ni) write_en_ff <= '0;
    else                       write_en_ff <= write_en_next;
  end
// END write_en

// START axil_if.bvalid
  logic bvalid_ff;
  logic bvalid_next;

  assign bvalid_next = write_state_next == StResp;

  always_ff @(posedge axil_if.clk_i or negedge axil_if.arst_ni) begin
    if      (!axil_if.arst_ni) bvalid_ff <= '0;
    else                       bvalid_ff <= bvalid_next;
  end
// END axil_if.bvalid

// START axil_if.awready
  logic awready_ff;
  logic awready_next;

  assign awready_next = read_state_next == StIdle;

  always_ff @(posedge axil_if.clk_i or negedge axil_if.arst_ni) begin
    if      (!axil_if.arst_ni) awready_ff <= '0;
    else                       awready_ff <= awready_next;
  end
// END axil_if.awready

// START data_out_ff
  axil_data_t data_out_ff;
  axil_data_t data_out_next;
  logic       data_out_en;

  assign      data_out_en   = write_state_next == StAddrData;
  assign      data_out_next = axil_if.wdata_i;

  always_ff @(posedge axil_if.clk_i or negedge axil_if.arst_ni) begin
    if      (!axil_if.arst_ni) data_out_ff <= '0;
    else if (data_out_en     ) data_out_ff <= data_out_next;
  end
// END data_ff

// START addr_write_ff
  native_addr_t addr_write_ff;
  native_addr_t addr_write_next;
  logic         addr_write_en;

  assign      addr_write_en   = write_state_next == StAddrData;
  assign      addr_write_next = axil2native_addr(axil_if.awaddr_i);

  always_ff @(posedge axil_if.clk_i or negedge axil_if.arst_ni) begin
    if      (!axil_if.arst_ni) addr_write_ff <= '0;
    else if (addr_write_en   ) addr_write_ff <= addr_write_next;
  end
// END addr_write_ff
// END write logic

// START out assignments
  assign native_if.addr_write   = addr_write_ff;
  assign native_if.addr_read    = addr_read_ff;
  assign native_if.read_en_sync = read_en_sync_ff;
  assign native_if.write_en     = write_en_ff;
  assign native_if.data2native  = data_out_ff;

  assign axil_if.arready_o = arready_ff;
  assign axil_if.awready_o = awready_ff;
  assign axil_if.wready_o  = awready_ff; // simultaneous with axil_if.awready
  assign axil_if.bvalid_o  = bvalid_ff;
  assign axil_if.rvalid_o  = rvalid_ff;
  assign axil_if.rdata_o   = rdata_ff;

  import vga_axil_pkg::axil_resp_t, vga_axil_pkg::OKAY;
  assign axil_if.rresp_o   = axil_resp_t'(OKAY);
  assign axil_if.bresp_o   = axil_resp_t'(OKAY);
// END out assignments

endmodule
