interface vga_arst_n_if (
  input logic clk
);
  logic arst_n;
endinterface
